// LA64 Privileged Instructions (Section 4.2)
// Note: All privileged instructions can ONLY be executed in PLV0

// 4.2.1 CSR访问指令 (use la64_csr_instr class)
`DEFINE_LA64_CSR_INSTR(CSRRD,   R2I14_TYPE, CSR, LA64, IMM)
`DEFINE_LA64_CSR_INSTR(CSRWR,   R2I14_TYPE, CSR, LA64, IMM)
`DEFINE_LA64_CSR_INSTR(CSRXCHG, R2I14_TYPE, CSR, LA64, IMM)

// 4.2.2 IOCSR访问指令 (use la64_privileged_instr class)
`DEFINE_LA64_PRIV_INSTR(IOCSRRD_B, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRRD_H, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRRD_W, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRRD_D, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRWR_B, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRWR_H, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRWR_W, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(IOCSRWR_D, R2_TYPE, SYSTEM, LA64)

// 4.2.3 Cache维护指令 (use la64_privileged_instr class)
`DEFINE_LA64_PRIV_INSTR(CACOP, R2I12_TYPE, SYSTEM, LA64, IMM)

// 4.2.4 TLB维护指令 (use la64_privileged_instr class)
`DEFINE_LA64_PRIV_INSTR(TLBSRCH,   R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(TLBRD,     R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(TLBWR,     R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(TLBFILL,   R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(TLBCLR,    R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(TLBFLUSH,  R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(INVTLB,    R3_TYPE, SYSTEM, LA64)

// 4.2.5 软件页表遍历指令 (use la64_privileged_instr class)
`DEFINE_LA64_PRIV_INSTR(LDDIR, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(LDPTE, R2_TYPE, SYSTEM, LA64)

// 4.2.6 其它杂项指令 (use la64_privileged_instr class)
`DEFINE_LA64_PRIV_INSTR(ERTN, R2_TYPE, SYSTEM, LA64)
`DEFINE_LA64_PRIV_INSTR(DBCL, R2_TYPE, SYSTEM, LA64, IMM)
`DEFINE_LA64_PRIV_INSTR(IDLE, R2_TYPE, SYSTEM, LA64, IMM)
