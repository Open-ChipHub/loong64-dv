// TODO: Add custom instruction name enum
