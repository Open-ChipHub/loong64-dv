//#########基础整数指令##########
// 加减法
`DEFINE_INSTR(ADD_W,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ADD_D,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(SUB_W,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(SUB_D,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ADDI_W, R2I12_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(ADDI_D, R2I12_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(ADDU16I_D, R2I16_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(ALSL_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ALSL_WU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ALSL_D, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(LU12I_W, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(LU32I_D, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(LU52I_D, R2I12_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(PCADDI, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(PCADDU12I, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(PCADDU18I, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(PCALAU12I, R1I21_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(NOP,    R2I12_TYPE, ARITHMETIC, LA64)
// 比较
`DEFINE_INSTR(SLT,      R3_TYPE, COMPARE, LA64)
`DEFINE_INSTR(SLTU,     R3_TYPE, COMPARE, LA64)
`DEFINE_INSTR(SLTI,  R2I12_TYPE, COMPARE, LA64, IMM)
`DEFINE_INSTR(SLTUI, R2I12_TYPE, COMPARE, LA64, IMM)
// 逻辑运算
`DEFINE_INSTR(AND,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(OR,      R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(NOR,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(XOR,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ANDN,    R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ORN,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ANDI, R2I12_TYPE, LOGICAL, LA64, UIMM)
`DEFINE_INSTR(ORI,  R2I12_TYPE, LOGICAL, LA64, UIMM)
`DEFINE_INSTR(XORI, R2I12_TYPE, LOGICAL, LA64, UIMM)

`DEFINE_INSTR(MUL_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MUL_D, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULH_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULH_WU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULH_D, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULH_DU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULW_D_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MULW_D_WU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(DIV_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(DIV_WU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(DIV_D, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(DIV_DU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MOD_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MOD_WU, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MOD_D, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MOD_DU, R3_TYPE, ARITHMETIC, LA64)
// 移位运算类指令
`DEFINE_INSTR(SLL_W, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SRL_W, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SRA_W, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(ROTR_W, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SLLI_W, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(SRLI_W, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(SRAI_W, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(ROTRI_W, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(SLL_D, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SRL_D, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SRA_D, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(ROTR_D, R3_TYPE, SHIFT, LA64)
`DEFINE_INSTR(SLLI_D, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(SRLI_D, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(SRAI_D, R2I12_TYPE, SHIFT, LA64, UIMM)
`DEFINE_INSTR(ROTRI_D, R2I12_TYPE, SHIFT, LA64, UIMM)
// 位操作指令
`DEFINE_INSTR(EXT_W_B, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(EXT_W_H, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CLO_W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CLO_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CLZ_W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CLZ_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CTO_W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CTO_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CTZ_W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(CTZ_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BYTEPICK_W, R3_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BYTEPICK_D, R3_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVB_2H, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVB_4H, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVB_2W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVB_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVH_2W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(REVH_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BITREV_4B, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BITREV_8B, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BITREV_W, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BITREV_D, R2_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(BSTRINS_W, R2I12_TYPE, BITOPERATION, LA64, UIMM)
`DEFINE_INSTR(BSTRINS_D, R2I12_TYPE, BITOPERATION, LA64, UIMM)
`DEFINE_INSTR(BSTRPICK_W, R2I12_TYPE, BITOPERATION, LA64, UIMM)
`DEFINE_INSTR(BSTRPICK_D, R2I12_TYPE, BITOPERATION, LA64, UIMM)
`DEFINE_INSTR(MASKEQZ, R3_TYPE, BITOPERATION, LA64)
`DEFINE_INSTR(MASKNEZ, R3_TYPE, BITOPERATION, LA64)
// 转移指令
`DEFINE_INSTR(BEQ,  R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BNE,  R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BLT,  R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BGE,  R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BLTU, R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BGEU, R2I16_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BEQZ, R1I21_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(BNEZ, R1I21_TYPE, BRANCH, LA64, IMM)
`DEFINE_INSTR(B,  I26_TYPE, JUMP, LA64, IMM)
`DEFINE_INSTR(BL, I26_TYPE, JUMP, LA64, IMM)
`DEFINE_INSTR(JIRL, R2I16_TYPE, JUMP, LA64, IMM)
// 普通访存指令
`DEFINE_INSTR(LD_B,  R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_BU, R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_H,  R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_HU, R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_W,  R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_WU, R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LD_D,  R2I12_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(ST_B,  R2I12_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(ST_H,  R2I12_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(ST_W,  R2I12_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(ST_D,  R2I12_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(LDX_B,  R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_BU, R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_H,  R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_HU, R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_W,  R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_WU, R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDX_D,  R3_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(STX_B,  R3_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(STX_H,  R3_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(STX_W,  R3_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(STX_D,  R3_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(LDPTR_W, R2I14_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(LDPTR_D, R2I14_TYPE, LOAD,  LA64, IMM)
`DEFINE_INSTR(STPTR_W, R2I14_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(STPTR_D, R2I14_TYPE, STORE, LA64, IMM)
`DEFINE_INSTR(PRELD,  R2I12_TYPE, LOAD, LA64, IMM)
`DEFINE_INSTR(PRELDX, R3_TYPE, LOAD, LA64, IMM)
