// 加减法
`DEFINE_INSTR(ADD_W,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ADD_D,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(SUB_W,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(SUB_D,     R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(ADDI_W, R2I12_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(ADDI_D, R2I12_TYPE, ARITHMETIC, LA64, IMM)
`DEFINE_INSTR(NOP,    R2I12_TYPE, ARITHMETIC, LA64)
// 比较
`DEFINE_INSTR(SLT,      R3_TYPE, COMPARE, LA64)
`DEFINE_INSTR(SLTU,     R3_TYPE, COMPARE, LA64)
`DEFINE_INSTR(SLTI,  R2I12_TYPE, COMPARE, LA64, IMM)
`DEFINE_INSTR(SLTUI, R2I12_TYPE, COMPARE, LA64, IMM)
// 逻辑运算
`DEFINE_INSTR(AND,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(OR,      R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(NOR,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(XOR,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ANDN,    R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ORN,     R3_TYPE, LOGICAL, LA64)
`DEFINE_INSTR(ANDI, R2I12_TYPE, LOGICAL, LA64, UIMM)
`DEFINE_INSTR(ORI,  R2I12_TYPE, LOGICAL, LA64, UIMM)
`DEFINE_INSTR(XORI, R2I12_TYPE, LOGICAL, LA64, UIMM)

`DEFINE_INSTR(MUL_W, R3_TYPE, ARITHMETIC, LA64)
`DEFINE_INSTR(MUL_D, R3_TYPE, ARITHMETIC, LA64)
