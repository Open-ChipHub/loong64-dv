/*
 * LoongArch 浮点指令定义
 */

// 浮点算术运算指令
`DEFINE_FP_INSTR(FADD_S, R3_TYPE, ARITHMETIC, LA64)
